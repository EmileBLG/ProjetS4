----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/17/2024 04:34:26 PM
-- Design Name: 
-- Module Name: package_LUT - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;


package package_LUT_actor is

    type P_LUT_MAP is array (natural range <>) of std_logic_vector (3 downto 0);
    type P_LUT_TILE is array (natural range <>) of std_logic_vector (3 downto 0);
    
    constant P_LUT_MAP_ACTOR_1 : P_LUT_MAP(0 to 4095) := ( --dessiner acteurs dans le coin en haut à gauche avec outil mathias
    --Liste des tuiles dans un acteur (le tuyau)
    (x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"8",x"8",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"7",x"7",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"7",x"7",x"7",x"7"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"7",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0"),(x"0",x"0",x"0",x"0",x"0",x"0",x"8",x"8",x"8",x"8",x"0",x"0",x"0",x"0",x"0",x"0")


    --Liste des tuiles dans un acteur (le flappy bird)
    (x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8"),(x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8"),(x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8"),(x"8",x"8",x"8",x"8",x"8",x"8",x"7",x"7",x"7",x"7",x"7",x"7",x"8",x"8",x"8",x"8"),(x"8",x"8",x"8",x"8",x"7",x"7",x"4",x"4",x"4",x"4",x"7",x"f",x"7",x"8",x"8",x"8"),(x"8",x"8",x"8",x"7",x"4",x"4",x"4",x"4",x"4",x"7",x"f",x"f",x"f",x"7",x"8",x"8"),(x"8",x"7",x"7",x"7",x"7",x"4",x"4",x"4",x"4",x"7",x"f",x"f",x"7",x"f",x"7",x"8"),(x"7",x"f",x"f",x"f",x"f",x"7",x"4",x"4",x"4",x"7",x"f",x"f",x"7",x"f",x"7",x"8"),(x"7",x"f",x"f",x"f",x"f",x"f",x"7",x"4",x"4",x"4",x"7",x"f",x"f",x"f",x"7",x"8"),(x"8",x"7",x"f",x"f",x"f",x"7",x"4",x"4",x"4",x"4",x"4",x"7",x"7",x"7",x"7",x"7"),(x"8",x"8",x"7",x"7",x"7",x"4",x"4",x"4",x"4",x"4",x"7",x"6",x"6",x"6",x"6",x"6"),(x"8",x"8",x"7",x"4",x"4",x"4",x"4",x"4",x"4",x"7",x"6",x"7",x"7",x"7",x"7",x"7"),(x"8",x"8",x"8",x"7",x"7",x"4",x"4",x"4",x"4",x"4",x"7",x"6",x"6",x"6",x"6",x"6"),(x"8",x"8",x"8",x"8",x"7",x"4",x"4",x"4",x"4",x"4",x"4",x"7",x"7",x"7",x"7",x"7"),(x"8",x"8",x"8",x"8",x"8",x"7",x"7",x"7",x"7",x"7",x"7",x"8",x"8",x"8",x"8",x"8"),(x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8",x"8")
    
    
    others => "0000"
    );
    
    constant P_LUT_TILE_ACTOR_1 : P_LUT_TILE(0 to 2047) := ( --liste des pixels dans une tuile


    
    others => "0000"
    );
    
    
    
end package package_LUT_actor;

------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;

package package_LUT_bg is

    type P_LUT_MAP_BG is array (natural range <>) of std_logic_vector (5 downto 0);
    constant P_LUT_MAP_BACKGROUND : P_LUT_MAP_BG(0 to 4095) := (

    --Ca c'est la composition de chaque tuile de background (8 tuiles total)
 --tile 0:
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"d",x"d"
 x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"d",x"d",x"d"
 
 x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 
 x"d",x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 
 x"d",x"4",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"4",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"4",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 
 
 --tile 1
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"f",x"f",x"d"
 x"d",x"d",x"d",x"f",x"f",x"d",x"d",x"d",x"d",x"d",x"f",x"f",x"f",x"f",x"f",x"d"
 x"d",x"d",x"c",x"f",x"f",x"f",x"f",x"c",x"c",x"c",x"f",x"f",x"f",x"f",x"f",x"d"
 x"d",x"d",x"c",x"d",x"f",x"f",x"f",x"d",x"d",x"c",x"c",x"f",x"f",x"f",x"d",x"d"
 
 x"f",x"f",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"f",x"f",x"f",x"f",x"c",x"d",x"c",x"c",x"d",x"d",x"c",x"c",x"c",x"c",x"d",x"d"
 x"f",x"f",x"f",x"f",x"c",x"c",x"c",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"f",x"f",x"f",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"c",x"d",x"d",x"d",x"d"
 
 x"f",x"f",x"c",x"c",x"d",x"d",x"d",x"c",x"c",x"d",x"d",x"c",x"c",x"c",x"d",x"d"
 x"d",x"c",x"c",x"c",x"c",x"c",x"c",x"d",x"d",x"d",x"c",x"c",x"c",x"c",x"d",x"d"
 x"d",x"c",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"c",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"c",x"c",x"c"
 
 x"d",x"d",x"c",x"c",x"c",x"c",x"c",x"c",x"c",x"d",x"d",x"d",x"c",x"c",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"c",x"c",x"c",x"c",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d",x"d"
 
 
 --tile 2
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"
 x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e",x"e"


 --tile 3
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4",x"4"
 
 
 --tile 4:
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b",x"b"
 
 
 --tile 5
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a"
 
 x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"8",x"a",x"a",x"a"
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a"
 
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a"
 x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a"
 x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a"
 
 x"a",x"a",x"a",x"a",x"8",x"8",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"a",x"a"
 x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"8",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"8"
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"8",x"8",x"8"
 x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a",x"a"
 
 
 --tile 6        
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 
 --tile 7        
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
 x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0",x"0"
    
    others => "000000"
    );
    
    type P_LUT_TILE_BG is array (natural range <>) of std_logic_vector (3 downto 0);
    constant P_LUT_TILE_BACKGROUND : P_LUT_TILE_BG(0 to 16383) := (

    --Ca c'est lees tuiles de background (e.g., tuile 1, tuile 2, tuile 3, etc., pour le background)
        "0001", "0001", "0001", "0001", "0001", "0011", "0011", "0001", "0001", "0011", "0011", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0011", "0011", "0001", "0011",
        "0011", "0011", "0011", "0011", "0001", "0001", "0011", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0011", "0011", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0011", "0011", "0011",
        "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0011", "0011", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0011",
        "0001", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0011", "0011", "0011", "0011", "0001", "0011", "0011", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0011",
        "0001", "0011", "0001", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
        
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0001", "0110", "0001", "0001", "0110", "0110",
        "0100", "0110", "0110", "0101", "0110", "0001", "0001", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0001", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0101", "0001", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0001", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0100", "0110", "0110",
        "0101", "0110", "0110", "0110", "0001", "0110", "0110", "0101", "0001", "0110", "0110", "0110", "0100", "0100", "0001", "0100",
        "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0100", "0110", "0110", "0110",
        "0110", "0110", "0001", "0110", "0100", "0001", "0110", "0110", "0110", "0001", "0100", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0100",
        "0110", "0101", "0001", "0110", "0110", "0001", "0001", "0110", "0110", "0110", "0101", "0110", "0101", "0001", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001",
        "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110",
        "0001", "0110", "0101", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0101", "0110", "0100", "0110",
        "0110", "0101", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0101", "0110", "0100", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0001", "0110", "0110",
        "0101", "0101", "0001", "0110", "0110", "0110", "0101", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001",
        "0001", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0001", "0110", "0110", "0001", "0110", "0110",
        
        "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0101", "0110", "0001", "0110",
        "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0101", "0110", "0110", "0001", "0110", "0110", "0101", "0110", "0110", "0100", "0001", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110",
        
        "0110", "0110", "0110", "0001", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0100",
        "0100", "0100", "0110", "0110", "0110", "0001", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110",
        "0110", "0110", "0101", "0110", "0110", "0110", "0101", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0100", "0110", "0100", "0110", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0100", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0100", "0101", "0110", "0110", "0001", "0110", "0100", "0110", "0110", "0101", "0110", "0110",
        "0110", "0110", "0001", "0110", "0110", "0110", "0001", "0001", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0101", "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110",
        
        "0110", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0001", "0001", "0101", "0110", "0110", "0110", "0001", "0001", "0110", "0001", "0001", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110",
        "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0001", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0001", "0101", "0110", "0110", "0001", "0110", "0110", "0001", "0110", "0001", "0001", "0001", "0110", "0110", "0110",
        "0110", "0001", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0101", "0001", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110",
        
        "0110", "0001", "0101", "0110", "0110", "0110", "0001", "0001", "0110", "0110", "0001", "0101", "0001", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0101", "0110", "0110", "0110", "0001", "0110",
        "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0100", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110",
        
        "0110", "0101", "0001", "0001", "0110", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0100", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0001", "0110", "0001", "0001", "0110", "0001", "0110",
        
        "0110", "0101", "0001", "0001", "0110", "0110", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0100", "0110", "0100", "0110", "0110", "0110", "0110", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0101", "0001", "0110",
        "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0001", "0110", "0110",
        
        "0110", "0101", "0001", "0001", "0110", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0101", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0001", "0001", "0110",
        
        "0110", "0101", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0001", "0110", "0110", "0001", "0101", "0110",
        "0110", "0100", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0101", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0001", "0110", "0001", "0110", "0110", "0110", "0001", "0110",
        
        "0110", "0001", "0101", "0001", "0110", "0001", "0001", "0110", "0001", "0110", "0001", "0110", "0110", "0001", "0100", "0101",
        "0110", "0001", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110",
        "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0110", "0001", "0001", "0110",
        
        "0110", "0001", "0101", "0001", "0110", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0001", "0100", "0001", "0001",
        "0110", "0110", "0100", "0101", "0110", "0100", "0001", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0100", "0110", "0001", "0001", "0110", "0110", "0001", "0001", "0110",
        
        "0110", "0110", "0001", "0101", "0110", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0100", "0001", "0110", "0110", "0110", "0100", "0110", "0110", "0101", "0110", "0001", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0001", "0110",
        
        "0110", "0001", "0001", "0101", "0110", "0001", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0100",
        "0100", "0001", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0100", "0001", "0110",
        
        "0110", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0001", "0110", "0101", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0100", "0110", "0110",
        
        "0110", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0101", "0001", "0110", "0001", "0001", "0110", "0001", "0001",
        "0001", "0110", "0110", "0110", "0100", "0101", "0100", "0110", "0100", "0110", "0110", "0110", "0110", "0101", "0110", "0100",
        "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0001", "0001", "0101", "0110", "0101", "0001", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0001", "0110",
        
        "0110", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0110", "0110", "0001", "0001", "0101", "0110", "0101",
        "0110", "0101", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0100", "0100", "0100", "0110", "0110", "0110", "0110",
        "0001", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0110", "0110", "0001", "0110", "0110", "0001", "0101", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0001",
        "0001", "0001", "0001", "0110", "0001", "0001", "0110", "0001", "0001", "0110", "0100", "0110", "0001", "0001", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0100", "0110", "0110", "0110",
        "0001", "0110", "0001", "0110", "0001", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0001", "0001", "0110", "0001", "0001", "0001",
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0100", "0110",
        "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110",
        "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0101", "0110", "0110", "0001", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0001", "0110", "0001", "0001",
        "0001", "0100", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0110", "0110", "0001", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0001", "0001", "0100", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0001", "0110", "0110", "0001", "0110", "0001", "0001", "0110", "0110", "0001", "0110", "0001", "0110", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0001", "0001", "0001", "0001", "0110",
        "0001", "0001", "0110", "0001", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0101", "0110", "0001", "0110", "0110",
        "0110", "0110", "0110", "0110", "0101", "0001", "0001", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0001", "0110", "0100", "0110", "0001", "0110", "0110", "0110", "0001", "0001", "0110", "0001", "0001", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0001",
        "0001", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0101", "0110", "0001", "0110",
        "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0001", "0110", "0001",
        "0110", "0001", "0001", "0110", "0001", "0110", "0100", "0110", "0001", "0001", "0001", "0110", "0110", "0110", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0001", "0001", "0001", "0110",
        "0001", "0001", "0110", "0001", "0110", "0110", "0110", "0110", "0001", "0110", "0001", "0001", "0110", "0101", "0001", "0001",
        "0001", "0001", "0100", "0001", "0001", "0001", "0110", "0001", "0001", "0001", "0110", "0110", "0001", "0110", "0100", "0110",
        "0001", "0100", "0110", "0110", "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0001", "0110",
        
        "0110", "0110", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0001",
        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0001", "0001", "0001", "0101", "0001",
        "0101", "0001", "0001", "0001", "0001", "0110", "0001", "0101", "0001", "0100", "0110", "0110", "0001", "0110", "0001", "0001",
        "0101", "0100", "0001", "0100", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0110", "0001", "0001", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0001", "0101", "0001", "0110", "0110", "0001", "0001", "0100", "0110", "0110", "0100", "0001", "0001", "0100", "0001",
        "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110",
        
    others => "0000"
    );
    
    
    
end package package_LUT_bg;

