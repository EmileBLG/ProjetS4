----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/17/2024 04:34:26 PM
-- Design Name: 
-- Module Name: package_LUT - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;


package package_LUT_actor is

    type P_LUT_MAP is array (natural range <>) of std_logic_vector (3 downto 0);
    type P_LUT_TILE is array (natural range <>) of std_logic_vector (3 downto 0);
    
    constant P_LUT_MAP_ACTOR_1 : P_LUT_MAP(0 to 4095) := (
    -- row 1 of 64
    --0                  4                    8                                         16                                        24                                  31  
    X"2",X"1",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    --32                                      40                                        48                                        56                                  63  
    X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    
    -- row 2 of 64
    --0                  4                    8                                         16                                        24                                  31  
    X"2",X"1",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    --32                                      40                                        48                                        56                                  63  
    X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    
    -- row 3 of 64
    --0                  4                    8                                         16                                        24                                  31  
    X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    --32                                      40                                        48                                        56                                  63  
    X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    
    others => "0000"
    );
    
    constant P_LUT_TILE_ACTOR_1 : P_LUT_TILE(0 to 2047) := (
    -- tile 0
    X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", X"0",X"0",X"0",X"0", 
    "0000","0001","1010","0011", "0100","0101","0110","0111", "0000","0001","1010","0011", "0100","0101","0110","0111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    -- tile 1
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    -- tile 2
    others => "0000"
    );
    
    
    
end package package_LUT_actor;

------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;

package package_LUT_bg is

    type P_LUT_MAP_BG is array (natural range <>) of std_logic_vector (5 downto 0);
    constant P_LUT_MAP_BACKGROUND : P_LUT_MAP_BG(0 to 4095) := (
    -- row 1 of 64
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    
    -- row 2 of 64
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    "000010","000001","000000","000011", "000100","000101","000110","001111", "000010","000001","000000","000011", "000100","000101","000110","001111",
    
    others => "000000"
    );
    
    type P_LUT_TILE_BG is array (natural range <>) of std_logic_vector (3 downto 0);
    constant P_LUT_TILE_BACKGROUND : P_LUT_TILE_BG(0 to 16383) := (
    -- tile 0
    "0000","0001","1010","0011", "0100","0101","0110","0111", "0000","0001","1010","0011", "0100","0101","0110","0111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    -- tile 1
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    "0000","0001","0010","0011", "0100","0101","0110","0111", "1000","1001","1010","1011", "1100","1101","1110","1111",
    
    -- tile 2
    others => "0000"
    );
    
    
    
end package package_LUT_bg;

